`ifdef __ICARUS__
    `ifndef INCLUDE_PARAMS
        `include "./src/def_params.v"
    `endif
`endif
`define DISPLAY(A) `ifdef SIMULATE $display("%0d\tMEMORY: ",$time,A); `endif

module memory(
    input wire clk,
    input wire reset,

    //interface pipeline in
    `ifdef SIMULATE
    input wire [`ADDR_SIZE : 0] PC_in,
    input wire [`INSTR_SIZE : 0] instr_in,
    `endif
    input wire [4:0] opcode_in,
    input wire [2:0] funct_in,
    input wire nop_instr_in,
    input wire [`EX_WIDTH : 0] exception_in,
    input wire exception_in_valid,
    input wire pipeline_in_valid,
    input wire [`REG_DATA_SIZE : 0] result_in,
    input wire [`ADDR_SIZE : 0] addr,
    input wire [`REG_ADDR_SIZE : 0] rd_addr_in,

    //Interface pipeline out
    `ifdef SIMULATE
    output reg [`ADDR_SIZE : 0] PC_out,
    output reg [`INSTR_SIZE : 0] instr_out,
    `endif
    output reg nop_instr_out,
    output reg [`REG_DATA_SIZE : 0] result_out,
    output reg [`REG_ADDR_SIZE : 0] rd_addr_out,
    output reg pipeline_out_valid,
    output reg [`EX_WIDTH : 0] exception_out,
    output reg exception_out_valid,

    //Interface dmem
    output reg [`ADDR_SIZE : 0] mem_addr,
    output reg [`INSTR_SIZE : 0 ] mem_wr_data,
    output reg mem_wr_enable,
    input wire [`INSTR_SIZE : 0 ] mem_rd_data,
    output reg mem_rd_enable,
    input wire mem_rd_ready,

    input wire flush,
    input wire stall_in,
    output reg stall_out
);

    reg [`EX_WIDTH : 0] exception_out_rg;
    reg exception_out_valid_rg;

    reg load_wait = 0;

    always@(*) begin
        if(pipeline_in_valid) begin
            mem_rd_enable = 0;
            mem_wr_enable = 1;
            load_wait = 0;
            stall_out = 0;
            if(exception_in_valid) begin
                exception_out_valid_rg = exception_in_valid;
                exception_out_rg = exception_in;
            end
            else if(opcode_in == `OP_LOAD) begin
                mem_addr = addr;
                mem_rd_enable = 1;
                load_wait = 1;
                stall_out = 1;
            end
            else if(opcode_in == `OP_STORE) begin
                mem_addr = addr;
                mem_wr_enable = 1;
            end
            else begin

            end
        end
    end

    always@(posedge(clk)) begin
        if(reset) begin
            pipeline_out_valid <= 0;
            `DISPLAY("Reset")
        end
        else if(flush) begin
            pipeline_out_valid <= 0;
            `DISPLAY("Flush")
        end
        else if(stall_in) begin
            pipeline_out_valid <= pipeline_out_valid;
            `DISPLAY("Stall")
        end
        else if(pipeline_in_valid) begin
            if(opcode_in == `OP_LOAD) begin
                if(load_wait == 1 && mem_rd_ready == 1) begin
                    result_out <= mem_rd_data;
                end
            end
            else begin
                result_out <= result_in;
            end
            advancePipeline;
            `ifdef SIMULATE 
            PC_out <= PC_in;
            instr_out <= instr_in;
            printDebug; 
            `endif
        end
    end

    task advancePipeline;
    begin
        pipeline_out_valid <= pipeline_in_valid;
        rd_addr_out <= rd_addr_in;
        nop_instr_out <= nop_instr_in;
        exception_out <= exception_out_rg;
        exception_out_valid <= exception_out_valid_rg;
    end
    endtask

`ifdef SIMULATE
    task printDebug;
    begin
        $strobe("%0d\t************MEMORY Firing************", $time);
        if(nop_instr_in)
            `DISPLAY("OP: NOP")
        else begin
            case (opcode_in)
                `OP_LOAD:   `DISPLAY("OP: LOAD")
                `OP_STORE:  `DISPLAY("OP: STORE")
                default:    `DISPLAY("OP: Unkown")
            endcase
        end
        $strobe("%0d\tMEMORY: PC: %h instr: %h", $time, PC_out, instr_out);
        $strobe("%0d\tMEMORY: Exception: %d(valid %b)", $time, exception_out, exception_out_valid);
    end
    endtask
`endif

endmodule // memory