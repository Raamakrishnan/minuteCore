`ifdef __ICARUS__
    `ifndef INCLUDE_PARAMS
        `include "./src/params.v"
    `endif
`endif

module imem(

);

endmodule // imem